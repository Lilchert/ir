`timescale 1ns / 1ps

module tb;
    // Тактовый сигнал и сброс
    reg rst = 1;
    reg clk = 0;

    // Сигналы управления
    reg valid = 0;
    reg [7:0] data = 8'h6D; // 'A' в ASCII

    // Выходные сигналы
    wire ready;
    wire uart_tx;

    wire [31:0] baudrate = 31'd9600;
    // Параметры тестирования
    localparam CLK_PERIOD = 40; // 25 МГц (40 нс)
    localparam BIT_TIME = 1000000000/9600; // 104166 нс для 9600 бод

    // Инициализация UART передатчика
    uart_tx uart_inst (
        .clk(clk),
        .rst(rst),
        .baudrate(baudrate),   // Тестируем на 9600 бод
        .data(data),
        .valid(valid),
        .parity_en(1'b1),  // Включена проверка чётности
        .parity_type(1'b1), // Чётная чётность
        .tx(uart_tx),
        .ready(ready)
    );

    // Генератор тактовой частоты
    always #(CLK_PERIOD/2) clk = ~clk;

    initial begin
        // Создание файла дампа для GTKWave
        $dumpfile("waves.vcd");
        $dumpvars(0, tb);

        // Последовательность тестирования
        $display("=== Начало теста UART передатчика ===");

        // Сброс
        #100 rst = 0;
        $display("[%0t] Сброс снят", $time);

        // Ожидание готовности
        wait(ready == 1);
        $display("[%0t] Устройство готово к передаче", $time);

        // Запуск передачи
        $display("[%0t] Начало передачи символа 'A' (0x41)", $time);
        valid = 1;
        #10; valid = 0;

        // Мониторинг состояния линии
        $display("Ожидаемая последовательность (LSB first):");
        $display("Старт(0) 1 0 0 0 0 0 1 0 Чётность(1) Стоп(1)");

        // Проверка старт-бита
        wait(uart_tx == 0);
        $display("[%0t] Старт-бит обнаружен", $time);

        // Проверка данных (LSB first)
        #(BIT_TIME*1.5); check_bit(0, 1); // Бит 0
        #BIT_TIME; check_bit(1, 0);       // Бит 1
        #BIT_TIME; check_bit(2, 0);       // Бит 2
        #BIT_TIME; check_bit(3, 0);       // Бит 3
        #BIT_TIME; check_bit(4, 0);       // Бит 4
        #BIT_TIME; check_bit(5, 0);       // Бит 5
        #BIT_TIME; check_bit(6, 1);       // Бит 6
        #BIT_TIME; check_bit(7, 0);       // Бит 7

        // Проверка бита чётности
        #BIT_TIME;
        if(uart_tx == 1'b1)
            $display("[%0t] Бит чётности корректен (1)", $time);
        else
            $error("Ошибка бита чётности!");

        // Проверка стоп-бита
        #BIT_TIME;
        if(uart_tx == 1'b1)
            $display("[%0t] Стоп-бит корректен", $time);
        else
            $error("Ошибка стоп-бита!");

        // Завершение
        #100000;
        $display("=== Тест завершён успешно ===");
        $finish;
    end

    // Задача для проверки битов
    task check_bit;
        input [2:0] bit_num;
        input expected;
        begin
            if(uart_tx === expected)
                $display("[%0t] Бит %0d: %b (корректно)", $time, bit_num, uart_tx);
            else
                $error("Бит %0d: ожидалось %b, получено %b", bit_num, expected, uart_tx);
        end
    endtask
endmodule
